VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 1500.000 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 1496.000 283.730 1500.000 ;
    END
  END CLK
  PIN OUT[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 779.320 1500.000 779.920 ;
    END
  END OUT[0]
  PIN OUT[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.850 1496.000 1176.130 1500.000 ;
    END
  END OUT[1]
  PIN OUT[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1460.130 0.000 1460.410 4.000 ;
    END
  END OUT[2]
  PIN OUT[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1379.080 1500.000 1379.680 ;
    END
  END OUT[3]
  PIN OUT[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 179.560 1500.000 180.160 ;
    END
  END OUT[4]
  PIN OUT[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END OUT[5]
  PIN OUT[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END OUT[6]
  PIN OUT[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.080 4.000 359.680 ;
    END
  END OUT[7]
  PIN OUT[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END OUT[8]
  PIN OUT[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 300.600 1500.000 301.200 ;
    END
  END OUT[9]
  PIN imem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1259.400 1500.000 1260.000 ;
    END
  END imem_data[0]
  PIN imem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END imem_data[10]
  PIN imem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1198.200 4.000 1198.800 ;
    END
  END imem_data[11]
  PIN imem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END imem_data[12]
  PIN imem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.090 1496.000 851.370 1500.000 ;
    END
  END imem_data[13]
  PIN imem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.210 0.000 1298.490 4.000 ;
    END
  END imem_data[14]
  PIN imem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.010 1496.000 1013.290 1500.000 ;
    END
  END imem_data[15]
  PIN imem_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 659.640 1500.000 660.240 ;
    END
  END imem_data[16]
  PIN imem_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 1496.000 770.410 1500.000 ;
    END
  END imem_data[17]
  PIN imem_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1319.240 4.000 1319.840 ;
    END
  END imem_data[18]
  PIN imem_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.410 0.000 1054.690 4.000 ;
    END
  END imem_data[19]
  PIN imem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.450 0.000 973.730 4.000 ;
    END
  END imem_data[1]
  PIN imem_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 839.160 4.000 839.760 ;
    END
  END imem_data[20]
  PIN imem_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 900.360 1500.000 900.960 ;
    END
  END imem_data[21]
  PIN imem_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 0.000 892.770 4.000 ;
    END
  END imem_data[22]
  PIN imem_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.890 1496.000 1095.170 1500.000 ;
    END
  END imem_data[23]
  PIN imem_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.370 0.000 1135.650 4.000 ;
    END
  END imem_data[24]
  PIN imem_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.170 0.000 1379.450 4.000 ;
    END
  END imem_data[25]
  PIN imem_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END imem_data[26]
  PIN imem_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 59.880 1500.000 60.480 ;
    END
  END imem_data[27]
  PIN imem_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1438.920 4.000 1439.520 ;
    END
  END imem_data[28]
  PIN imem_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 958.840 4.000 959.440 ;
    END
  END imem_data[29]
  PIN imem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END imem_data[2]
  PIN imem_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 1496.000 201.850 1500.000 ;
    END
  END imem_data[30]
  PIN imem_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END imem_data[31]
  PIN imem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.810 1496.000 1257.090 1500.000 ;
    END
  END imem_data[3]
  PIN imem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.330 1496.000 526.610 1500.000 ;
    END
  END imem_data[4]
  PIN imem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1139.720 1500.000 1140.320 ;
    END
  END imem_data[5]
  PIN imem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.050 1496.000 932.330 1500.000 ;
    END
  END imem_data[6]
  PIN imem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 1496.000 39.930 1500.000 ;
    END
  END imem_data[7]
  PIN imem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END imem_data[8]
  PIN imem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 1496.000 364.690 1500.000 ;
    END
  END imem_data[9]
  PIN init_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1499.690 1496.000 1499.970 1500.000 ;
    END
  END init_addr[0]
  PIN init_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 0.000 487.050 4.000 ;
    END
  END init_addr[1]
  PIN init_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 1020.040 1500.000 1020.640 ;
    END
  END init_addr[2]
  PIN init_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.330 0.000 1216.610 4.000 ;
    END
  END init_addr[3]
  PIN init_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 1496.000 689.450 1500.000 ;
    END
  END init_addr[4]
  PIN init_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 420.280 1500.000 420.880 ;
    END
  END init_addr[5]
  PIN init_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END init_addr[6]
  PIN init_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END init_addr[7]
  PIN init_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1078.520 4.000 1079.120 ;
    END
  END init_en
  PIN mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END mem_addr[0]
  PIN mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END mem_addr[1]
  PIN mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.730 1496.000 1419.010 1500.000 ;
    END
  END mem_addr[2]
  PIN mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.770 1496.000 1338.050 1500.000 ;
    END
  END mem_addr[3]
  PIN mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 1496.000 445.650 1500.000 ;
    END
  END mem_addr[4]
  PIN mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.290 1496.000 607.570 1500.000 ;
    END
  END mem_addr[5]
  PIN mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 0.000 810.890 4.000 ;
    END
  END mem_addr[6]
  PIN mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END mem_addr[7]
  PIN mem_wr
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 1496.000 120.890 1500.000 ;
    END
  END mem_wr
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1496.000 539.960 1500.000 540.560 ;
    END
  END reset
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1488.080 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1488.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1488.080 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1494.080 1487.925 ;
      LAYER met1 ;
        RECT 0.070 10.240 1499.990 1488.480 ;
      LAYER met2 ;
        RECT 0.100 1495.720 39.370 1496.000 ;
        RECT 40.210 1495.720 120.330 1496.000 ;
        RECT 121.170 1495.720 201.290 1496.000 ;
        RECT 202.130 1495.720 283.170 1496.000 ;
        RECT 284.010 1495.720 364.130 1496.000 ;
        RECT 364.970 1495.720 445.090 1496.000 ;
        RECT 445.930 1495.720 526.050 1496.000 ;
        RECT 526.890 1495.720 607.010 1496.000 ;
        RECT 607.850 1495.720 688.890 1496.000 ;
        RECT 689.730 1495.720 769.850 1496.000 ;
        RECT 770.690 1495.720 850.810 1496.000 ;
        RECT 851.650 1495.720 931.770 1496.000 ;
        RECT 932.610 1495.720 1012.730 1496.000 ;
        RECT 1013.570 1495.720 1094.610 1496.000 ;
        RECT 1095.450 1495.720 1175.570 1496.000 ;
        RECT 1176.410 1495.720 1256.530 1496.000 ;
        RECT 1257.370 1495.720 1337.490 1496.000 ;
        RECT 1338.330 1495.720 1418.450 1496.000 ;
        RECT 1419.290 1495.720 1499.410 1496.000 ;
        RECT 0.100 4.280 1499.960 1495.720 ;
        RECT 0.650 4.000 80.770 4.280 ;
        RECT 81.610 4.000 161.730 4.280 ;
        RECT 162.570 4.000 242.690 4.280 ;
        RECT 243.530 4.000 323.650 4.280 ;
        RECT 324.490 4.000 404.610 4.280 ;
        RECT 405.450 4.000 486.490 4.280 ;
        RECT 487.330 4.000 567.450 4.280 ;
        RECT 568.290 4.000 648.410 4.280 ;
        RECT 649.250 4.000 729.370 4.280 ;
        RECT 730.210 4.000 810.330 4.280 ;
        RECT 811.170 4.000 892.210 4.280 ;
        RECT 893.050 4.000 973.170 4.280 ;
        RECT 974.010 4.000 1054.130 4.280 ;
        RECT 1054.970 4.000 1135.090 4.280 ;
        RECT 1135.930 4.000 1216.050 4.280 ;
        RECT 1216.890 4.000 1297.930 4.280 ;
        RECT 1298.770 4.000 1378.890 4.280 ;
        RECT 1379.730 4.000 1459.850 4.280 ;
        RECT 1460.690 4.000 1499.960 4.280 ;
      LAYER met3 ;
        RECT 4.000 1439.920 1496.000 1488.005 ;
        RECT 4.400 1438.520 1496.000 1439.920 ;
        RECT 4.000 1380.080 1496.000 1438.520 ;
        RECT 4.000 1378.680 1495.600 1380.080 ;
        RECT 4.000 1320.240 1496.000 1378.680 ;
        RECT 4.400 1318.840 1496.000 1320.240 ;
        RECT 4.000 1260.400 1496.000 1318.840 ;
        RECT 4.000 1259.000 1495.600 1260.400 ;
        RECT 4.000 1199.200 1496.000 1259.000 ;
        RECT 4.400 1197.800 1496.000 1199.200 ;
        RECT 4.000 1140.720 1496.000 1197.800 ;
        RECT 4.000 1139.320 1495.600 1140.720 ;
        RECT 4.000 1079.520 1496.000 1139.320 ;
        RECT 4.400 1078.120 1496.000 1079.520 ;
        RECT 4.000 1021.040 1496.000 1078.120 ;
        RECT 4.000 1019.640 1495.600 1021.040 ;
        RECT 4.000 959.840 1496.000 1019.640 ;
        RECT 4.400 958.440 1496.000 959.840 ;
        RECT 4.000 901.360 1496.000 958.440 ;
        RECT 4.000 899.960 1495.600 901.360 ;
        RECT 4.000 840.160 1496.000 899.960 ;
        RECT 4.400 838.760 1496.000 840.160 ;
        RECT 4.000 780.320 1496.000 838.760 ;
        RECT 4.000 778.920 1495.600 780.320 ;
        RECT 4.000 720.480 1496.000 778.920 ;
        RECT 4.400 719.080 1496.000 720.480 ;
        RECT 4.000 660.640 1496.000 719.080 ;
        RECT 4.000 659.240 1495.600 660.640 ;
        RECT 4.000 599.440 1496.000 659.240 ;
        RECT 4.400 598.040 1496.000 599.440 ;
        RECT 4.000 540.960 1496.000 598.040 ;
        RECT 4.000 539.560 1495.600 540.960 ;
        RECT 4.000 479.760 1496.000 539.560 ;
        RECT 4.400 478.360 1496.000 479.760 ;
        RECT 4.000 421.280 1496.000 478.360 ;
        RECT 4.000 419.880 1495.600 421.280 ;
        RECT 4.000 360.080 1496.000 419.880 ;
        RECT 4.400 358.680 1496.000 360.080 ;
        RECT 4.000 301.600 1496.000 358.680 ;
        RECT 4.000 300.200 1495.600 301.600 ;
        RECT 4.000 240.400 1496.000 300.200 ;
        RECT 4.400 239.000 1496.000 240.400 ;
        RECT 4.000 180.560 1496.000 239.000 ;
        RECT 4.000 179.160 1495.600 180.560 ;
        RECT 4.000 120.720 1496.000 179.160 ;
        RECT 4.400 119.320 1496.000 120.720 ;
        RECT 4.000 60.880 1496.000 119.320 ;
        RECT 4.000 59.480 1495.600 60.880 ;
        RECT 4.000 10.715 1496.000 59.480 ;
      LAYER met4 ;
        RECT 602.895 13.095 635.040 1167.385 ;
        RECT 637.440 13.095 711.840 1167.385 ;
        RECT 714.240 13.095 788.640 1167.385 ;
        RECT 791.040 13.095 865.440 1167.385 ;
        RECT 867.840 13.095 942.240 1167.385 ;
        RECT 944.640 13.095 1019.040 1167.385 ;
        RECT 1021.440 13.095 1095.840 1167.385 ;
        RECT 1098.240 13.095 1110.145 1167.385 ;
  END
END user_proj_example
END LIBRARY

