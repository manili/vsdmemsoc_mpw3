magic
tech sky130A
magscale 1 2
timestamp 1636138118
<< obsli1 >>
rect 1104 2159 298816 297585
<< obsm1 >>
rect 14 2048 299998 297696
<< metal2 >>
rect 7930 299200 7986 300000
rect 24122 299200 24178 300000
rect 40314 299200 40370 300000
rect 56690 299200 56746 300000
rect 72882 299200 72938 300000
rect 89074 299200 89130 300000
rect 105266 299200 105322 300000
rect 121458 299200 121514 300000
rect 137834 299200 137890 300000
rect 154026 299200 154082 300000
rect 170218 299200 170274 300000
rect 186410 299200 186466 300000
rect 202602 299200 202658 300000
rect 218978 299200 219034 300000
rect 235170 299200 235226 300000
rect 251362 299200 251418 300000
rect 267554 299200 267610 300000
rect 283746 299200 283802 300000
rect 299938 299200 299994 300000
rect 18 0 74 800
rect 16210 0 16266 800
rect 32402 0 32458 800
rect 48594 0 48650 800
rect 64786 0 64842 800
rect 80978 0 81034 800
rect 97354 0 97410 800
rect 113546 0 113602 800
rect 129738 0 129794 800
rect 145930 0 145986 800
rect 162122 0 162178 800
rect 178498 0 178554 800
rect 194690 0 194746 800
rect 210882 0 210938 800
rect 227074 0 227130 800
rect 243266 0 243322 800
rect 259642 0 259698 800
rect 275834 0 275890 800
rect 292026 0 292082 800
<< obsm2 >>
rect 20 299144 7874 299200
rect 8042 299144 24066 299200
rect 24234 299144 40258 299200
rect 40426 299144 56634 299200
rect 56802 299144 72826 299200
rect 72994 299144 89018 299200
rect 89186 299144 105210 299200
rect 105378 299144 121402 299200
rect 121570 299144 137778 299200
rect 137946 299144 153970 299200
rect 154138 299144 170162 299200
rect 170330 299144 186354 299200
rect 186522 299144 202546 299200
rect 202714 299144 218922 299200
rect 219090 299144 235114 299200
rect 235282 299144 251306 299200
rect 251474 299144 267498 299200
rect 267666 299144 283690 299200
rect 283858 299144 299882 299200
rect 20 856 299992 299144
rect 130 800 16154 856
rect 16322 800 32346 856
rect 32514 800 48538 856
rect 48706 800 64730 856
rect 64898 800 80922 856
rect 81090 800 97298 856
rect 97466 800 113490 856
rect 113658 800 129682 856
rect 129850 800 145874 856
rect 146042 800 162066 856
rect 162234 800 178442 856
rect 178610 800 194634 856
rect 194802 800 210826 856
rect 210994 800 227018 856
rect 227186 800 243210 856
rect 243378 800 259586 856
rect 259754 800 275778 856
rect 275946 800 291970 856
rect 292138 800 299992 856
<< metal3 >>
rect 0 287784 800 287904
rect 299200 275816 300000 275936
rect 0 263848 800 263968
rect 299200 251880 300000 252000
rect 0 239640 800 239760
rect 299200 227944 300000 228064
rect 0 215704 800 215824
rect 299200 204008 300000 204128
rect 0 191768 800 191888
rect 299200 180072 300000 180192
rect 0 167832 800 167952
rect 299200 155864 300000 155984
rect 0 143896 800 144016
rect 299200 131928 300000 132048
rect 0 119688 800 119808
rect 299200 107992 300000 108112
rect 0 95752 800 95872
rect 299200 84056 300000 84176
rect 0 71816 800 71936
rect 299200 60120 300000 60240
rect 0 47880 800 48000
rect 299200 35912 300000 36032
rect 0 23944 800 24064
rect 299200 11976 300000 12096
<< obsm3 >>
rect 800 287984 299200 297601
rect 880 287704 299200 287984
rect 800 276016 299200 287704
rect 800 275736 299120 276016
rect 800 264048 299200 275736
rect 880 263768 299200 264048
rect 800 252080 299200 263768
rect 800 251800 299120 252080
rect 800 239840 299200 251800
rect 880 239560 299200 239840
rect 800 228144 299200 239560
rect 800 227864 299120 228144
rect 800 215904 299200 227864
rect 880 215624 299200 215904
rect 800 204208 299200 215624
rect 800 203928 299120 204208
rect 800 191968 299200 203928
rect 880 191688 299200 191968
rect 800 180272 299200 191688
rect 800 179992 299120 180272
rect 800 168032 299200 179992
rect 880 167752 299200 168032
rect 800 156064 299200 167752
rect 800 155784 299120 156064
rect 800 144096 299200 155784
rect 880 143816 299200 144096
rect 800 132128 299200 143816
rect 800 131848 299120 132128
rect 800 119888 299200 131848
rect 880 119608 299200 119888
rect 800 108192 299200 119608
rect 800 107912 299120 108192
rect 800 95952 299200 107912
rect 880 95672 299200 95952
rect 800 84256 299200 95672
rect 800 83976 299120 84256
rect 800 72016 299200 83976
rect 880 71736 299200 72016
rect 800 60320 299200 71736
rect 800 60040 299120 60320
rect 800 48080 299200 60040
rect 880 47800 299200 48080
rect 800 36112 299200 47800
rect 800 35832 299120 36112
rect 800 24144 299200 35832
rect 880 23864 299200 24144
rect 800 12176 299200 23864
rect 800 11896 299120 12176
rect 800 2143 299200 11896
<< metal4 >>
rect 4208 2128 4528 297616
rect 19568 2128 19888 297616
rect 34928 2128 35248 297616
rect 50288 2128 50608 297616
rect 65648 2128 65968 297616
rect 81008 2128 81328 297616
rect 96368 2128 96688 297616
rect 111728 2128 112048 297616
rect 127088 2128 127408 297616
rect 142448 2128 142768 297616
rect 157808 2128 158128 297616
rect 173168 2128 173488 297616
rect 188528 2128 188848 297616
rect 203888 2128 204208 297616
rect 219248 2128 219568 297616
rect 234608 2128 234928 297616
rect 249968 2128 250288 297616
rect 265328 2128 265648 297616
rect 280688 2128 281008 297616
rect 296048 2128 296368 297616
<< obsm4 >>
rect 120579 2619 127008 233477
rect 127488 2619 142368 233477
rect 142848 2619 157728 233477
rect 158208 2619 173088 233477
rect 173568 2619 188448 233477
rect 188928 2619 203808 233477
rect 204288 2619 219168 233477
rect 219648 2619 222029 233477
<< labels >>
rlabel metal2 s 56690 299200 56746 300000 6 CLK
port 1 nsew signal input
rlabel metal3 s 299200 155864 300000 155984 6 OUT[0]
port 2 nsew signal output
rlabel metal2 s 235170 299200 235226 300000 6 OUT[1]
port 3 nsew signal output
rlabel metal2 s 292026 0 292082 800 6 OUT[2]
port 4 nsew signal output
rlabel metal3 s 299200 275816 300000 275936 6 OUT[3]
port 5 nsew signal output
rlabel metal3 s 299200 35912 300000 36032 6 OUT[4]
port 6 nsew signal output
rlabel metal3 s 0 95752 800 95872 6 OUT[5]
port 7 nsew signal output
rlabel metal2 s 64786 0 64842 800 6 OUT[6]
port 8 nsew signal output
rlabel metal3 s 0 71816 800 71936 6 OUT[7]
port 9 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 OUT[8]
port 10 nsew signal output
rlabel metal3 s 299200 60120 300000 60240 6 OUT[9]
port 11 nsew signal output
rlabel metal3 s 299200 251880 300000 252000 6 imem_data[0]
port 12 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 imem_data[10]
port 13 nsew signal input
rlabel metal3 s 0 239640 800 239760 6 imem_data[11]
port 14 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 imem_data[12]
port 15 nsew signal input
rlabel metal2 s 170218 299200 170274 300000 6 imem_data[13]
port 16 nsew signal input
rlabel metal2 s 259642 0 259698 800 6 imem_data[14]
port 17 nsew signal input
rlabel metal2 s 202602 299200 202658 300000 6 imem_data[15]
port 18 nsew signal input
rlabel metal3 s 299200 131928 300000 132048 6 imem_data[16]
port 19 nsew signal input
rlabel metal2 s 154026 299200 154082 300000 6 imem_data[17]
port 20 nsew signal input
rlabel metal3 s 0 263848 800 263968 6 imem_data[18]
port 21 nsew signal input
rlabel metal2 s 210882 0 210938 800 6 imem_data[19]
port 22 nsew signal input
rlabel metal2 s 194690 0 194746 800 6 imem_data[1]
port 23 nsew signal input
rlabel metal3 s 0 167832 800 167952 6 imem_data[20]
port 24 nsew signal input
rlabel metal3 s 299200 180072 300000 180192 6 imem_data[21]
port 25 nsew signal input
rlabel metal2 s 178498 0 178554 800 6 imem_data[22]
port 26 nsew signal input
rlabel metal2 s 218978 299200 219034 300000 6 imem_data[23]
port 27 nsew signal input
rlabel metal2 s 227074 0 227130 800 6 imem_data[24]
port 28 nsew signal input
rlabel metal2 s 275834 0 275890 800 6 imem_data[25]
port 29 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 imem_data[26]
port 30 nsew signal input
rlabel metal3 s 299200 11976 300000 12096 6 imem_data[27]
port 31 nsew signal input
rlabel metal3 s 0 287784 800 287904 6 imem_data[28]
port 32 nsew signal input
rlabel metal3 s 0 191768 800 191888 6 imem_data[29]
port 33 nsew signal input
rlabel metal3 s 0 143896 800 144016 6 imem_data[2]
port 34 nsew signal input
rlabel metal2 s 40314 299200 40370 300000 6 imem_data[30]
port 35 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 imem_data[31]
port 36 nsew signal input
rlabel metal2 s 251362 299200 251418 300000 6 imem_data[3]
port 37 nsew signal input
rlabel metal2 s 105266 299200 105322 300000 6 imem_data[4]
port 38 nsew signal input
rlabel metal3 s 299200 227944 300000 228064 6 imem_data[5]
port 39 nsew signal input
rlabel metal2 s 186410 299200 186466 300000 6 imem_data[6]
port 40 nsew signal input
rlabel metal2 s 7930 299200 7986 300000 6 imem_data[7]
port 41 nsew signal input
rlabel metal2 s 18 0 74 800 6 imem_data[8]
port 42 nsew signal input
rlabel metal2 s 72882 299200 72938 300000 6 imem_data[9]
port 43 nsew signal input
rlabel metal2 s 299938 299200 299994 300000 6 init_addr[0]
port 44 nsew signal input
rlabel metal2 s 97354 0 97410 800 6 init_addr[1]
port 45 nsew signal input
rlabel metal3 s 299200 204008 300000 204128 6 init_addr[2]
port 46 nsew signal input
rlabel metal2 s 243266 0 243322 800 6 init_addr[3]
port 47 nsew signal input
rlabel metal2 s 137834 299200 137890 300000 6 init_addr[4]
port 48 nsew signal input
rlabel metal3 s 299200 84056 300000 84176 6 init_addr[5]
port 49 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 init_addr[6]
port 50 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 init_addr[7]
port 51 nsew signal input
rlabel metal3 s 0 215704 800 215824 6 init_en
port 52 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 mem_addr[0]
port 53 nsew signal output
rlabel metal2 s 129738 0 129794 800 6 mem_addr[1]
port 54 nsew signal output
rlabel metal2 s 283746 299200 283802 300000 6 mem_addr[2]
port 55 nsew signal output
rlabel metal2 s 267554 299200 267610 300000 6 mem_addr[3]
port 56 nsew signal output
rlabel metal2 s 89074 299200 89130 300000 6 mem_addr[4]
port 57 nsew signal output
rlabel metal2 s 121458 299200 121514 300000 6 mem_addr[5]
port 58 nsew signal output
rlabel metal2 s 162122 0 162178 800 6 mem_addr[6]
port 59 nsew signal output
rlabel metal3 s 0 119688 800 119808 6 mem_addr[7]
port 60 nsew signal output
rlabel metal2 s 24122 299200 24178 300000 6 mem_wr
port 61 nsew signal output
rlabel metal3 s 299200 107992 300000 108112 6 reset
port 62 nsew signal input
rlabel metal4 s 4208 2128 4528 297616 6 vccd1
port 63 nsew power input
rlabel metal4 s 34928 2128 35248 297616 6 vccd1
port 63 nsew power input
rlabel metal4 s 65648 2128 65968 297616 6 vccd1
port 63 nsew power input
rlabel metal4 s 96368 2128 96688 297616 6 vccd1
port 63 nsew power input
rlabel metal4 s 127088 2128 127408 297616 6 vccd1
port 63 nsew power input
rlabel metal4 s 157808 2128 158128 297616 6 vccd1
port 63 nsew power input
rlabel metal4 s 188528 2128 188848 297616 6 vccd1
port 63 nsew power input
rlabel metal4 s 219248 2128 219568 297616 6 vccd1
port 63 nsew power input
rlabel metal4 s 249968 2128 250288 297616 6 vccd1
port 63 nsew power input
rlabel metal4 s 280688 2128 281008 297616 6 vccd1
port 63 nsew power input
rlabel metal4 s 19568 2128 19888 297616 6 vssd1
port 64 nsew ground input
rlabel metal4 s 50288 2128 50608 297616 6 vssd1
port 64 nsew ground input
rlabel metal4 s 81008 2128 81328 297616 6 vssd1
port 64 nsew ground input
rlabel metal4 s 111728 2128 112048 297616 6 vssd1
port 64 nsew ground input
rlabel metal4 s 142448 2128 142768 297616 6 vssd1
port 64 nsew ground input
rlabel metal4 s 173168 2128 173488 297616 6 vssd1
port 64 nsew ground input
rlabel metal4 s 203888 2128 204208 297616 6 vssd1
port 64 nsew ground input
rlabel metal4 s 234608 2128 234928 297616 6 vssd1
port 64 nsew ground input
rlabel metal4 s 265328 2128 265648 297616 6 vssd1
port 64 nsew ground input
rlabel metal4 s 296048 2128 296368 297616 6 vssd1
port 64 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 300000 300000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 66858312
string GDS_START 938140
<< end >>

